package Testbench;

import UART::*;  
import StmtFSM::*;


module mkTb(Empty);
    

endmodule: mkTb





endpackage: Testbench